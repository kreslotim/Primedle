    Mac OS X            	   2  �     �                                    ATTR;���  �   �   s                  �   9  com.apple.quarantine   )     com.apple.lastuseddate#PS 7D-  9   *  $com.apple.metadata:_kMDItemUserTags F0083;623322c1;Safari;D6E03F4D-8DB5-417D-8AD6-FBFB36815F45!8Tb    �el    bplist00�                            	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            This resource fork intentionally left blank                                                                                                                                                                                                                            ��