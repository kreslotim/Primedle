    Mac OS X            	   2  �     �                                    ATTR;���  �   �   �                  �   9  com.apple.quarantine        com.apple.lastuseddate#PS 57-  %   H  com.apple.macl 7E0083;623c964d;Safari;E00B97E3-2F48-4857-BD4B-2173528413E5�<Tb    ��     �"2�aL���s���;�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        This resource fork intentionally left blank                                                                                                                                                                                                                            ��