    Mac OS X            	   2  �     �                                    ATTR;���  �   �   s                  �   9  com.apple.quarantine   )     com.apple.lastuseddate#PS 05-  9   *  $com.apple.metadata:_kMDItemUserTags 40083;62332086;Safari;1359B7D1-776F-4005-813B-4A4666A6E2DAߧ8b    �})    bplist00�                            	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            This resource fork intentionally left blank                                                                                                                                                                                                                            ��