    Mac OS X            	   2  �     �                                    ATTR;���  �   �   I                  �   9  com.apple.quarantine    �     com.apple.lastuseddate#PS 57-0083;623c964d;Safari;E00B97E3-2F48-4857-BD4B-2173528413E5a:Tb    �P�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          This resource fork intentionally left blank                                                                                                                                                                                                                            ��